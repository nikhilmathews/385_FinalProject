/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  maze_RAM
(
		input [9:0] read_addressX, read_addressY, Pac_X_Pos, Pac_Y_Pos, Ghost_X_Pos, Ghost_Y_Pos,
		output logic data_Out, up_wall, down_wall, left_wall ,right_wall, up_wall_g, down_wall_g , left_wall_g, right_wall_g
);

// mem has width of 3 bits and a total of 400 addresses
logic [479:0][639:0] mem = {
640'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
640'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
640'b 0000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000,
640'b 0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000,
640'b 0000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000,
640'b 0000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000,
640'b 0000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000,
640'b 0000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000,
640'b 0000001111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111000000,
640'b 0000111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111110000,
640'b 0000111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011111000000000000001111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111110000000000111110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110111110000000000000000000000000000000000000000000000000011111011111111111111111111111111111111111111111111111111111111111111111111111110111110000000000000000000000000000000000000000000000000011111011111101111100000000000000000000000000000000000000000000000000111110111111111111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000000000111110111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000001111100000000000111111000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000001111110000000000011111000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011110000,
640'b 0000111110000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000111110000,
640'b 0000001111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000000000000000000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111000000,
640'b 0000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000000000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000,
640'b 0000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000,
640'b 0000000111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110000000,
640'b 0000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000,
640'b 0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000,
640'b 0000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000,
640'b 0000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000011111100000000000011111100000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111101111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111011111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
640'b 0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
640'b 0000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000001111100000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000011111000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111110000000000111110000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000111110000000000111110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110000000000000000000000000000000000000000000000000011111011111101111100000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000011111011111101111100000000000000000000000000000000000000000000000000111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000,
640'b 0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
640'b 0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000,
640'b 0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
640'b 0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000001111100000000000111111000000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000001111110000000000011111000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000,
640'b 0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000,
640'b 0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
640'b 0000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000,
640'b 0000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000,
640'b 0000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000,
640'b 0000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000,
640'b 0000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000011111100000000000011111000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000001111100000000000011111100000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000,
640'b 0000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000,
640'b 0000000111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011110000000,
640'b 0000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000,
640'b 0000011111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111100000,
640'b 0000111100000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000011110000,
640'b 0000111100000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111000000000000001111100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111110000000000111110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000011110000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000111100000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000011110000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111100000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000011110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000111100000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000011110000,
640'b 0000111100000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000011110000,
640'b 0000111100000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000011110000,
640'b 0000111100000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000011110000,
640'b 0000111100000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000001111100000000000011111000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000001111100000000000011111000000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000001111100000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000011111000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000011111000000000001111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111000000000001111100000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000001111100000000011110000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000111100000000011111000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000,
640'b 0000111100000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000011110000,
640'b 0000111100000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000011110000,
640'b 0000111100000000111110111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111110111110000000000000000000000111110111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110111110000000011110000,
640'b 0000111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000,
640'b 0000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000011101111011110100111111101111011101101111010011111100101111111110011101101110111110100011111011110100111110000000000000000000000111110001010111111111101111101110111010111101101011111111111100000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000011111101100011110011101111111011111010101101001100001000111110000000000000000000000111110011111010110011111111110011111101110001111001101111001111011111110111111111110110001011010011111111100000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000001111100000000000011111000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011110000,
640'b 0000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011110000,
640'b 0000111100000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000011110000,
640'b 0000111100000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000011110000,
640'b 0000011111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111100000,
640'b 0000000111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000,
640'b 0000000111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011110000000,
640'b 0000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000,
640'b 0000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000,
640'b 0000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000,
640'b 0000000000001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000,
640'b 0000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000,
};

//initial
//begin
//
////	 $readmemb("sprite_bytes/maze.txt", mem);
//end


parameter [9:0] pac_size = 10'd18;
parameter [9:0] Ghost_size = 10'd18;
parameter [9:0] mid = 10'd9;
always_comb
 begin
	data_Out<= mem[read_addressY][read_addressX];
	if (Pac_Y_Pos > 10'd0)
		up_wall <= mem[Pac_Y_Pos-10'd02][Pac_X_Pos] | mem[Pac_Y_Pos-10'd02][Pac_X_Pos + mid] | mem[Pac_Y_Pos-10'd02][Pac_X_Pos + pac_size] ;
	else 
		up_wall <= 1'b1;
	if (Pac_Y_Pos < (10'd479 - pac_size))
		down_wall <= mem[Pac_Y_Pos+10'd02+pac_size][Pac_X_Pos] | mem[Pac_Y_Pos+10'd02+pac_size][Pac_X_Pos + mid] | mem[Pac_Y_Pos+10'd02+pac_size][Pac_X_Pos + pac_size];
	else 
		down_wall <= 1'b1;
	if (Pac_X_Pos > 10'd0)
		left_wall <= mem[Pac_Y_Pos][Pac_X_Pos-10'd02] | mem[Pac_Y_Pos + mid][Pac_X_Pos-10'd02] | mem[Pac_Y_Pos + pac_size][Pac_X_Pos-10'd02] ;
	else 
		left_wall <= 1'b1;
	if (Pac_X_Pos < (10'd639 - pac_size))
		right_wall <= mem[Pac_Y_Pos][Pac_X_Pos+10'd02+pac_size] | mem[Pac_Y_Pos + mid][Pac_X_Pos+10'd02+pac_size] | mem[Pac_Y_Pos + pac_size][Pac_X_Pos+10'd02+pac_size];
	else 
		right_wall <= 1'b1;	

	if (Ghost_Y_Pos > 10'd0)
		up_wall_g <= mem[Ghost_Y_Pos-10'd02][Ghost_X_Pos]| mem[Ghost_Y_Pos-10'd02][Ghost_X_Pos + mid] | mem[Ghost_Y_Pos-10'd02][Ghost_X_Pos + pac_size] ;
	else 
		up_wall_g <= 1'b1;
	if (Ghost_Y_Pos < (10'd479 - Ghost_size))
		down_wall_g <= mem[Ghost_Y_Pos+10'd02+Ghost_size][Ghost_X_Pos] | mem[Ghost_Y_Pos+10'd02+pac_size][Ghost_X_Pos + mid] | mem[Ghost_Y_Pos+10'd02+pac_size][Ghost_X_Pos + pac_size];
	else 
		down_wall_g <= 1'b1;
	if (Ghost_X_Pos > 10'd0)
		left_wall_g <= mem[Ghost_Y_Pos][Ghost_X_Pos-10'd02]  | mem[Ghost_Y_Pos + mid][Ghost_X_Pos-10'd02] | mem[Ghost_Y_Pos + pac_size][Ghost_X_Pos-10'd02] ;
	else 
		left_wall_g <= 1'b1;
	if (Ghost_X_Pos < (10'd639 - Ghost_size))
		right_wall_g <= mem[Ghost_Y_Pos][Ghost_X_Pos+10'd02+Ghost_size] | mem[Ghost_Y_Pos + mid][Ghost_X_Pos+10'd02+pac_size] | mem[Ghost_Y_Pos + pac_size][Ghost_X_Pos+10'd02+pac_size];
	else 
		right_wall_g <= 1'b1;	

end


endmodule
